module tb;
    initial begin
        $display("Hello World! Icarus Verilog is working.");
        $finish; // This ends the simulation
    end
endmodule